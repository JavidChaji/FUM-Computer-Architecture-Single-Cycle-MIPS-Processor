//memory unit
module IMemBank(input memread, input [15:0] address, output reg [15:0] readdata);
 
  reg [15:0] mem_array [255:0];
  
//   integer i;
  initial begin
     /* mem_array[0] = 16'b0000000001010000;		// $2 = $0 + $1
		mem_array[1] = 16'b0001000011001010;		// $3 = $0 + 10
		mem_array[2] = 16'b0001011011000101;		// $3 = $3 + 5
		mem_array[3] = 16'b1000000100000000;		// $4 = mem 0($0) 
		mem_array[4] = 16'b1001000001100100;		// beq $0, $1, -4
		mem_array[5] = 16'b1111000000000000;		// jump 0;*/
				//			algoritm test
	/*	mem_array[0] = 16'b0001001001001010;		// addi $1, $1, 10
		mem_array[1] = 16'b0001001010010100;		// addi $2, $1, 20
		mem_array[2] = 16'b0000001010011000;		//	add $3, $1, $2
		mem_array[3] = 16'b1000000011000000;		// mem 0($0) = $3
		mem_array[4] = 16'b0111000001000000;		// $1 = mem 0($0)
		mem_array[5] = 16'b0001001101001010;		// addi $5, $1, 10;
		mem_array[6] = 16'b0000001010100010;		// and $4, $1, $2
		mem_array[7] = 16'b0000001010101011;		// or $5, $1, $2
		mem_array[8] = 16'b0000001010110100;		//	xor $6, $1, $2
		mem_array[9] = 16'b0000001010111101;		// xnor $7, $1, $2
		mem_array[10] = 16'b0000001010100110;		// slt $4, $1, $2
		mem_array[11] = 16'b0010001101111111;		// andi $5, $1, 63
		mem_array[12] = 16'b0011001110000000;		// ori $6, $1, 0
		mem_array[13] = 16'b0100001111001010;		// subi $7, $1, 10
		mem_array[14] = 16'b1111000000000000;		// jump 0		*/
		
		
		/* A[10];									mod
			for(int i=0; i<6; i++)
				A[i] = 2;
			for(int i=6; i<10; i++)
				A[i] = 1;
			for(int i=0; i<10; i++)
				for(int j=i+1; i<10; j++){
					if(A[j]<A[i]){
						int temp = A[j];
						A[j] = A[i];
						A[i] = temp;
					}
				}
				
			int x = 1, maxX = 1, mod = A[0];
			for(int i=0; i<9; i++){
				if(A[i+1]==A[i])
					x++;
				else{
					if(x > maxX){
						maxX = x;
						mod = A[i];
						}
					x = 1;
				}
			}
			
			if(x > maxX){
						maxX = x;
						mod = A[i];
				}
			*/
							
						// A -> $7										algoritm mod
			/*mem_array[0] = 16'b0001000001000000;	//	addi $1, $0, 0			
			mem_array[1] = 16'b0001000010000101;	// addi $2, $0, 5
			mem_array[2] = 16'b0001000011000010;	// addi $3, $0, 2
			mem_array[3] = 16'b1100001010000100;	// bgt $1, $2, 4
			mem_array[4] = 16'b0000001111100000;	// add $4, $1, $7
			mem_array[5] = 16'b1000100011000000;	//	sw $3, 0($4)
			mem_array[6] = 16'b0001001001000001; 	// addi $1, $1, 1;
			mem_array[7] = 16'b1111000000000011; 	// jump 3;
			
			mem_array[8] = 16'b0001000001000110;	//	addi $1, $0, 6
			mem_array[9] = 16'b0001000010001001;	// addi $2, $0, 9
			mem_array[10] = 16'b0001000011000001;	// addi $3, $0, 1
			mem_array[11] = 16'b1100001010000100;	// bgt $1, $2, 4
			mem_array[12] = 16'b0000001111100000;	// add $4, $1, $7
			mem_array[13] = 16'b1000100011000000;	//	sw $3, 0($4)
			mem_array[14] = 16'b0001001001000001; 	// addi $1, $1, 1;
			mem_array[15] = 16'b1111000000001011; 	// jump 11;
			
			mem_array[16] = 16'b0001000001000000;	//	addi $1, $0, 0
			mem_array[17] = 16'b0001000010001001;	// addi $2, $0, 9
			mem_array[18] = 16'b1100001010010001;	// bgt $1, $2, 17
			mem_array[19] = 16'b0001001101000001; 	// addi $5, $1, 1
			mem_array[20] = 16'b1100101010001101;	// bgt $5, $2, 13
			mem_array[21] = 16'b0000001111011000; 	// add $3, $1, $7		A[i]
			mem_array[22] = 16'b0000101111100000;	// add $4, $5, $7
			mem_array[23] = 16'b0111011011000000;	// lw $3 ,0($3)
			mem_array[24] = 16'b0111100100000000; 	// lw $4, 0($4)
			mem_array[25] = 16'b0001011011111111;	// addi $3, $3, -1
			mem_array[26] = 16'b1100100011000101;	// bgt $4, $3, 5
			mem_array[27] = 16'b0001011110000000;	// addi $6, $3, 0
			mem_array[28] = 16'b0000001111011000;	//	addi $3, $1, $7
			mem_array[29] = 16'b1000011100000000;	// sw $4, 0($3)
			mem_array[30] = 16'b0000101111100000;	// add $4, $5, $7
			mem_array[31] = 16'b1000100110000000;	// sw $6, 0($4)
			mem_array[32] = 16'b0001101101000001;	// addi $5, $5, 1;
			mem_array[33] = 16'b1111000000010100;	// jump 20
			mem_array[34] = 16'b0001001001000001; 	// addi $1, $1, 1
			mem_array[35] = 16'b1111000000010010;	// jump 18
			
			mem_array[36] = 16'b0001000010000001; 	//	addi $2, $0, 1
			mem_array[37] = 16'b0001000011000001;	// addi $3, $0, 1
			mem_array[38] = 16'b0001000001000000; 	// addi $1, $0, 0;
			mem_array[39] = 16'b0001000100001000;	// addi $4, $0, 8;
			mem_array[40] = 16'b1100001100001111;	//	bgt $1, $4, 15
			mem_array[41] = 16'b0000001111101000;	// add $5, $1, $7
			mem_array[42] = 16'b0111101101000000;	// lw $5, 0($5)
			mem_array[43] = 16'b0001001110000001;	// addi $6, $1, 1;
			mem_array[44] = 16'b0000110111110000;	//	add $6, $6, $7
			mem_array[45] = 16'b0111110110000000;	// lw $6, 0($6)
			mem_array[46] = 16'b1010101110000010;	// bnq $5, $6, 2
			mem_array[47] = 16'b0001010010000001;	// addi $2, $2, 1
			mem_array[48] = 16'b1111000000110110;	// jump 54
			mem_array[49] = 16'b1100011010000010;	// bgt $3, $2, 2
			mem_array[50] = 16'b0000010000011000;	// add $3, $2, $0
			mem_array[51] = 16'b0000000101100000;	// add $4, $0, $5
			mem_array[52] = 16'b0001000010000001;	// addi $2 , $0, 1
			mem_array[53] = 16'b0001000100001000;	// addi $4, $0, 8;
			mem_array[54] = 16'b0001001001000001;	// addi $1, $1, 1
			mem_array[55] = 16'b1111000000101000;	// jump 40	
			
			mem_array[56] = 16'b1100011010000010;	// bgt $3, $2, 2
			mem_array[57] = 16'b0000010000011000;	// add $3, $2, $0
			mem_array[58] = 16'b0000000101100000;	// add $4, $0, $5	*/
			
			/* 
				for(int i=0; i<10; i++)
					A[i] = i;
				int max = A[0], min=A[0]
				for(int i=0; i<10; i++){
					if(A[i] > max)
						max = A[i];
					if(A[i] < min)
						min = A[i];
				}
			*/
					// A -> $7				algoritm max, min
			// mem_array[0] = 16'b0001_000_001_000000;		// addi $1, $0, 0
			// mem_array[1] = 16'b0001_000_110_001001;		//	addi $6, $0, 9
			// mem_array[2] = 16'b1100_001_110_000100;		//	bgt $1, $6, 4
			// mem_array[3] = 16'b0000_001_111_010_000;		//	add $2, $1, $7
			// mem_array[4] = 16'b1000_010_001_000000;		//	sw $1, 0($2)
			// mem_array[5] = 16'b0001_001_001_000001;		//	addi $1, $1, 1
			// mem_array[6] = 16'b1111_000000000010;		// jump 2
		
			// mem_array[7] = 16'b0111_111011000000;		// lw $3, 0($7) 
			// mem_array[8] = 16'b0111_111100000000;		//	lw $4, 0($7)
			// mem_array[9] = 16'b0001_000001000000;		//	addi $1, $0, 0
			// mem_array[10] = 16'b1100_001110001000;		//	bgt $1, $6, 8
			// mem_array[11] = 16'b0000_001111010000;		//	add	$2, $1, $7
			// mem_array[12] = 16'b0111_010101000000;		//	lw $5, 0($2)
			// mem_array[13] = 16'b1011_101011000001;		//	blt $5, $3, 1 
			// mem_array[14] = 16'b0001_101011000000;		//	addi $3, $5, 0
			// mem_array[15] = 16'b1100_101100000001;		//	bgt $5, $4, 1 
			// mem_array[16] = 16'b0001_101100000000;		// addi $4, $5, 0
			// mem_array[17] = 16'b0001_001001000001;		// addi $1, $1, 1
			// mem_array[18] = 16'b1111_000000001010;		// jump 10

			// mem_array[19] = 16'b0000_011000011000;		// add $3, $3, $0
			// mem_array[20] = 16'b0000_100000100000;		// add $4, $4, $0


		// int n = 8;
		// int max=0;
		// int min=16'b1111_1111_1111_1111;
		// for(int i = 0 ; i <= n;i++){
		//     if(ar[i] > max){
		//         max = ar[i];
		//     }
		//     if(ar[i] < min){
		//         min = ar[i];
		//     }
		// }



		// i = $1
		// n = $6
		// min = $3
		// max = $4
		// temp1 = $2
		// temp2 = $5
		// baseReg = $7

		mem_array[0] <= 16'b0001_000_001_000000;// addi $1, $0, 0
		mem_array[1] <= 16'b0001_000_110_001000;// addi $6, $0, 8

		mem_array[2]  <= 16'b0001_000_001_000000;// addi $1, $0, 0

		mem_array[3] <= 16'b0001_000_100_000000;// addi $4, $0, 0
		mem_array[4] <= 16'b0010_000_111_000000;// andi $7, $0, 0
		mem_array[5] <= 16'b0001_000_011_011111;// addi $3, $0, 65535 but 63

		mem_array[6] <= 16'b1100_001_110_001000;// bgt $1, $6, 8
		mem_array[7] <= 16'b0000_111_001_010_000;// add $2, $7, $1
		mem_array[8] <= 16'b0111_010_101_000000;// lhw $5, 0($2)

		mem_array[9] <= 16'b1011_101_100_000001;// blt $5, $4, 1
		mem_array[10] <= 16'b0000_000_101_100_000;// add $4, $0 ,$5 

		mem_array[11] <= 16'b1100_101_011_000001;// bgt $5, $3, 1
		mem_array[12] <= 16'b0000_000_101_011_000;// add $3, $0, $5

		mem_array[13] <= 16'b0001_001_001_000001;// addi $1, $1, 1

		mem_array[14] <= 16'b1111_000000000110;// jump 5

		mem_array[15] <= 16'b0001_000_010_010011;// addi $2, $0, 19
		mem_array[16] <= 16'b0001_000_101_010100;// addi $5, $0, 20

		mem_array[17] <= 16'b1000_010_011_000000;// shw $3, 0($2)
		mem_array[18] <= 16'b1000_101_100_000000;// shw $4, 0($5)





		mem_array[19] <= 16'b0011_011_111_000111;// ori $7, $3, 7 //ori check
		mem_array[20] <= 16'b0100_111_010_000001;// subi $2, $7, 1 //subi check
		mem_array[21] <= 16'b1001_100_011_000010;// beq $4, $3,2   //beq check
		mem_array[22] <= 16'b0001_000_000_000000;// addi $0, $0, 0
		mem_array[23] <= 16'b0001_011_011_000001;// addi $3, $3, 1
		mem_array[24] <= 16'b1010_100_011_111100;// bne $4, $3, -4 //bne check
	


	end
 
  always@(memread, address, mem_array[address])
  begin
    if(memread)begin
      readdata=mem_array[address];
    end
  end

endmodule
