module ALU(input [15:0] data1,data2,input [3:0] aluoperation,output reg [15:0] result,output reg zero,lt,gt);

  always@(*)
  begin
    case (aluoperation)
      4'b0000 : result = data1 + data2; // ADD
      4'b0001 : result = data1 - data2; // SUB
      4'b0010 : result = data1 & data2; // AND
      4'b0011 : result = data1 | data2; // OR
      4'b0100 : result = data1 ^ data2; // XOR
		  4'b0101 : result = ~(data1 ^ data2); //XNOR
		  4'b0110 : result = data1<data2 ? 16'b1 : 16'b0;	// slt
      default : result = data1 + data2; // ADD
    endcase
    
    if(data1>data2)
		begin
		 zero = 1'b0;
       gt = 1'b1;
       lt = 1'b0; 
      end else if(data1<data2)
      begin
		 zero = 1'b0;
       gt = 1'b0;
       lt = 1'b1;  
      end
      else 
		begin
			zero = 1'b1;
			gt = 1'b0;
			lt = 1'b0;
		end
     
  end
  

endmodule
